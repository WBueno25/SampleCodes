/*/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
 ////////////////////////////////////////////////// LOGIC UNIT ////////////////////////////////////////////////////////////////
 //////////////////////////////////////// Developed By: Willian Analdo Nunes ///////////////////////////////////////////////////
 //////////////////////////////////////////// PUCRS, Porto Alegre, 2020      ///////////////////////////////////////////////////
 /////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////*/

`include "pkg.sv"
import my_pkg::*;

module logicUnit
    (input logic clk,
    input logic [31:0]  opA,
    input logic [31:0]  opB,
    input               instruction_type i,
    output logic [31:0] result_out);

    logic [31:0]        result;

    always_comb
        if(i==OP0)             // XOR 
            result <= opA ^ opB;
        else if(i==OP1)         // OR 
            result <= opA | opB;
        else                   // AND
            result <= opA & opB;

    always @(posedge clk)
        result_out <= result;

endmodule
