/*/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
 ////////////////////////////////////////////////// BYPASS UNIT ////////////////////////////////////////////////////////////////
 //////////////////////////////////////// Developed By: Willian Analdo Nunes ///////////////////////////////////////////////////
 //////////////////////////////////////////// PUCRS, Porto Alegre, 2020      ///////////////////////////////////////////////////
 /////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////*/

`include "pkg.sv"
import my_pkg::*;

module bypassUnit                   // LUI, NOP E INVALID
    (input logic clk,
    input logic reset,
    input logic [31:0]  opA,
    output logic [31:0] result_out);

    always @(posedge clk or negedge reset)
        if(!reset)
            result_out <= '0;
        else
            result_out <= opA;

endmodule